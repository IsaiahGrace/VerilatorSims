
typedef logic [7:0] word;
typedef logic [4:0] address;
              
