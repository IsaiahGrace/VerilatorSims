
typedef logic [7:0] word;
